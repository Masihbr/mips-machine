module control();
endmodule