module EXE_to_MEM();

endmodule

        .mem_write(mem_write_MEM),
        .alu_result(alu_result_MEM),
        .is_LB_SB(is_LB_SB_MEM),
        .rt_data(rt_data_MEM),
        .mem_data_out(mem_data_out_MEM),
        .cache_en(cache_en_MEM),
        .clk(clk),
        .rst_b(rst_b)